LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TWO_COMP IS PORT
(
  A : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
  A_COMP: OUT STD_LOGIC_VECTOR(64 DOWNTO 0)
);
END ENTITY TWO_COMP;

ARCHITECTURE BEHAVIORAL OF TWO_COMP IS
SIGNAL A_NOT, A_COMP_TEMP: STD_LOGIC_VECTOR(63 DOWNTO 0);
BEGIN
  A_NOT <= NOT(A);
  A_COMP_TEMP <= STD_LOGIC_VECTOR(SIGNED(A_NOT) + 1);
  A_COMP <= STD_LOGIC_VECTOR(RESIZE(SIGNED(A_COMP_TEMP), A_COMP'LENGTH));
END BEHAVIORAL;
