LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY HALF_ADDER IS PORT
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END ENTITY HALF_ADDER;

ARCHITECTURE BEHAVIORAL OF HALF_ADDER IS 
BEGIN
  S <= A XOR B;
  C <= A AND B;
END BEHAVIORAL;
