LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RC_ADDER_64 IS PORT
(
  A,B: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
  S  : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END ENTITY RC_ADDER_64;

ARCHITECTURE BEHAVIORAL OF RC_ADDER_64 IS
SIGNAL A_TEMP, B_TEMP, C_TEMP, S_TEMP: STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS => '0');

COMPONENT HALF_ADDER PORT
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END COMPONENT;
  
COMPONENT FULL_ADDER PORT
(
  A,B,CI: IN STD_LOGIC;
  S, CO: OUT STD_LOGIC
);
END COMPONENT;

BEGIN
  A_TEMP <= A;
  B_TEMP <= B;

  -- FIRT INPUT IS HALF ADDER
  HA_0: HALF_ADDER PORT MAP
    (
      A  => A_TEMP(0),
      B  => B_TEMP(0),
      S  => S_TEMP(0),
      C  => C_TEMP(0)
    );

  -- SUBSEQUENT FULL ADDER CHAIN
  FA_CHAIN: FOR I IN 1 TO 63 GENERATE
    FA_I: FULL_ADDER PORT MAP
      (
	A  => A_TEMP(I),
   	B  => B_TEMP(I),
	CI => C_TEMP(I-1),
	S  => S_TEMP(I),
	CO => C_TEMP(I)
      );
  END GENERATE FA_CHAIN;

  -- ASSIGNING OUTPUT
  S <= S_TEMP;
END BEHAVIORAL;