LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY COMPRESSOR_ADDER IS
GENERIC
(
  INPUT_WIDTH: INTEGER := 64
);
PORT 
(
  Cin       : IN STD_LOGIC;
  V, W, X, Y: IN STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0);
  Cout      : OUT STD_LOGIC;
  SUM       : OUT STD_LOGIC_VECTOR(INPUT_WIDTH DOWNTO 0)
);
END ENTITY COMPRESSOR_ADDER;

ARCHITECTURE BEHAVIORAL OF COMPRESSOR_ADDER IS
SIGNAL Cin_TEMP, RCA_C_TEMP: STD_LOGIC := '0';
SIGNAL V_TEMP, W_TEMP, X_TEMP, Y_TEMP, C_TEMP, S_TEMP: STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
SIGNAL Cout_TEMP, SUM_TEMP: STD_LOGIC_VECTOR(INPUT_WIDTH DOWNTO 0):= (OTHERS => '0') ;

COMPONENT RIPPLE_CARRY_ADDER PORT 
(
  A,B  : IN STD_LOGIC_VECTOR(62 DOWNTO 0);
  S    : OUT STD_LOGIC_VECTOR(62 DOWNTO 0);
  CARRY: OUT STD_LOGIC
);
END COMPONENT;

COMPONENT COMPRESSOR PORT
(
  V, W, X, Y, Cin: IN STD_LOGIC;
  Cout, C, S     : OUT STD_LOGIC
);
END COMPONENT;

COMPONENT FULL_ADDER PORT
(
  A,B,CI: IN STD_LOGIC;
  S, CO : OUT STD_LOGIC
);
END COMPONENT;

BEGIN

 -- ASSIGN INPUTS
 Cin_TEMP <= Cin;
 V_TEMP   <= V;
 W_TEMP   <= W;
 X_TEMP   <= X;
 Y_TEMP   <= Y;

 -- LAYER 0: COMPRESSORS LAYER
 COMP_0: COMPRESSOR PORT MAP
   (
     V    => V_TEMP(0),
	 W    => W_TEMP(0),
	 X    => X_TEMP(0),
	 Y    => Y_TEMP(0),
	 Cin  => Cin_TEMP,
	 Cout => Cout_TEMP(0),
	 C    => C_TEMP(0),
	 S    => S_TEMP(0)
   );
	 
 COMPRESSOR_LAYER: FOR I IN 1 TO INPUT_WIDTH-1 GENERATE
   COMP_I: COMPRESSOR PORT MAP 
    (
	  V    => V_TEMP(I),
	  W    => W_TEMP(I),
	  X    => X_TEMP(I),
	  Y    => Y_TEMP(I),
	  Cin  => Cout_TEMP(I-1),
	  Cout => Cout_TEMP(I),
	  C    => C_TEMP(I),
	  S    => S_TEMP(I)
	);
  END GENERATE;

  -- RIPPLE CARRY ADDER LAYER
  SUM_TEMP(0) <= S_TEMP(0);
  
  RCA: RIPPLE_CARRY_ADDER PORT MAP
   (
     A     => S_TEMP(INPUT_WIDTH-1 DOWNTO 1),
	 B     => C_TEMP(INPUT_WIDTH-2 DOWNTO 0),
	 S     => SUM_TEMP(INPUT_WIDTH-1 DOWNTO 1),
	 CARRY => RCA_C_TEMP
	);
	
  -- ONE FINAL ADDER TO ADD ALL THE CARRY TERMS OF LAST BLOCK
  FA: FULL_ADDER PORT MAP
   (
     A  => RCA_C_TEMP,
	 B  => C_TEMP(INPUT_WIDTH-1),
	 CI => C_TEMP(INPUT_WIDTH-1),
	 S  => SUM_TEMP(INPUT_WIDTH),
	 CO => Cout_TEMP(INPUT_WIDTH)
	);
	
  -- ASSIGNING OUTPUT
  SUM  <= SUM_TEMP;
  Cout <= Cout_TEMP(INPUT_WIDTH);
  
END BEHAVIORAL;
	 