LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CS_ADDER IS
GENERIC
(
  INPUT_WIDTH : INTEGER := 64
);

PORT
(
  X,Y,Z : IN STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0);
  S     : OUT STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0);
  CO    : OUT STD_LOGIC
);
END ENTITY CS_ADDER;

ARCHITECTURE BEHAVIORAL OF CS_ADDER IS
SIGNAL X_TEMP, Y_TEMP, Z_TEMP, 
S0_TEMP, C0_TEMP: STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0):= (OTHERS => '0');

SIGNAL S1_TEMP, C1_TEMP: STD_LOGIC_VECTOR(INPUT_WIDTH DOWNTO 0) := (OTHERS => '0');

COMPONENT FULL_ADDER PORT
(
  A,B,CI: IN STD_LOGIC;
  S, CO: OUT STD_LOGIC
);
END COMPONENT;

COMPONENT HALF_ADDER PORT
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END COMPONENT;

BEGIN
  X_TEMP <= X;
  Y_TEMP <= Y;
  Z_TEMP <= Z;

  -- CHAIN OF FULL ADDERS TO PRODUCE C AND S
  CSA_CHAIN: FOR I IN 0 TO INPUT_WIDTH-1 GENERATE
    FA_I: FULL_ADDER PORT MAP
      (
	A  => X_TEMP(I),
	B  => Y_TEMP(I),
	CI => Z_TEMP(I),
	S  => S0_TEMP(I),
	CO => C0_TEMP(I)
      );
  END GENERATE CSA_CHAIN;

  -- RIPPLE CARRY SECTION
  S1_TEMP(0) <= S0_TEMP(0);
  C1_TEMP(0) <= C0_TEMP(0);

  -- FIRST NODE WITH HALF ADDER
  HA_1: HALF_ADDER PORT MAP
    (
      A => C0_TEMP(0),
      B => S0_TEMP(1),
      S => S1_TEMP(1),
      C => C1_TEMP(1)
    );

  RC_FULL_ADDERS: FOR I IN 2 TO INPUT_WIDTH-1 GENERATE
   FA_I: FULL_ADDER PORT MAP
     (
       A  => C0_TEMP(I-1),
       B  => S0_TEMP(I),
       CI => C1_TEMP(I-1),
       S  => S1_TEMP(I),
       CO => C1_TEMP(I)
     );
   END GENERATE RC_FULL_ADDERS;

  -- LAST STAGE CARRY HALF ADDER
  HA_64: HALF_ADDER PORT MAP
    (
      A => C0_TEMP(63),
      B => C1_TEMP(63),
      S => S1_TEMP(64),
      C => C1_TEMP(64)
    );

  -- ASSIGINING OUTPUT
  S  <= S1_TEMP(INPUT_WIDTH-1 DOWNTO 0);
  CO <= C1_TEMP(64);
    
END BEHAVIORAL;
