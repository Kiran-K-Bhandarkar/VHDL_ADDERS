LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HC_ADDER IS
GENERIC
(
  INPUT_WIDTH : INTEGER := 64
);

PORT
(
  A,B : IN STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0);
  S   : OUT STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0)
);
END ENTITY HC_ADDER;

ARCHITECTURE BEHAVIORAL OF HC_ADDER IS
SIGNAL A_TEMP, B_TEMP, S_TEMP,
P0_TEMP, G0_TEMP, P1_TEMP, G1_TEMP,
P2_TEMP, G2_TEMP, P3_TEMP, G3_TEMP,
P4_TEMP, G4_TEMP, P5_TEMP, G5_TEMP,
P6_TEMP, G6_TEMP, P7_TEMP, G7_TEMP: STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0):= (OTHERS => '0');

COMPONENT HALF_ADDER PORT 
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END COMPONENT;

COMPONENT PROCESS_ELEMENT PORT
(
  Gi, Gj, Pi, Pj: IN STD_LOGIC;
  P, G: OUT STD_LOGIC
);
END COMPONENT;

BEGIN
  A_TEMP <= A;
  B_TEMP <= B;

  -- STAGE 0: OUTPUT FROM THE HALF ADDERS - PREPOCESSING STAGE
  PRE_PROCESSING: FOR I IN 0 TO INPUT_WIDTH-1 GENERATE
    HA_I: HALF_ADDER PORT MAP 
	(
	  A => A_TEMP(I), B => B_TEMP(I), 
	  S => P0_TEMP(I), C => G0_TEMP(I)
	);
  END GENERATE PRE_PROCESSING;

  -- STAGE 1
  P1_TEMP(0) <= P0_TEMP(0);
  G1_TEMP(0) <= G0_TEMP(0);

  -- NODE 2,4,6....62
  EVEN_NODES_S1: FOR I IN 1 TO (INPUT_WIDTH/2)-1 GENERATE
    P1_TEMP(2*I) <= P0_TEMP(2*I);
    G1_TEMP(2*I) <= G0_TEMP(2*I);
  END GENERATE EVEN_NODES_S1;

  -- NODE 3,5,7....63
  ODD_NODES_S1: FOR I IN 0 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S1_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G0_TEMP((2*I)+1),
	Pi => P0_TEMP((2*I)+1),
	Gj => G0_TEMP((2*I)),
	Pj => P0_TEMP((2*I)),
	P  => P1_TEMP((2*I)+1),
	G  => G1_TEMP((2*I)+1)
      );
   END GENERATE ODD_NODES_S1;

  -- STAGE 2
  -- NODE 0,1,2
  STAGE_2_INIT: FOR I IN 0 TO 2 GENERATE
    P2_TEMP(I) <= P1_TEMP(I);
    G2_TEMP(I) <= G1_TEMP(I);
  END GENERATE STAGE_2_INIT;

  -- NODE 4,6,8....62
  EVEN_NODES_S2: FOR I IN 2 TO (INPUT_WIDTH/2)-1 GENERATE
    P2_TEMP(2*I) <= P1_TEMP(2*I);
    G2_TEMP(2*I) <= G1_TEMP(2*I);
  END GENERATE EVEN_NODES_S2;

  -- NODE 3,5,7....63
  ODD_NODES_S2: FOR I IN 1 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S2_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G1_TEMP((2*I)+1),
	Pi => P1_TEMP((2*I)+1),
	Gj => G1_TEMP((2*I)-1),
	Pj => P1_TEMP((2*I)-1),
	P  => P2_TEMP((2*I)+1),
	G  => G2_TEMP((2*I)+1)
      );
   END GENERATE ODD_NODES_S2;

  -- STAGE 3
  -- NODE 0,1,2....4
  STAGE_3_INIT: FOR I IN 0 TO 4 GENERATE
    P3_TEMP(I) <= P2_TEMP(I);
    G3_TEMP(I) <= G2_TEMP(I);
  END GENERATE STAGE_3_INIT;
  
  -- NODE 6,8,10...62
  EVEN_NODES_S3: FOR I IN 3 TO (INPUT_WIDTH/2)-1 GENERATE
    P3_TEMP(2*I) <= P2_TEMP(2*I);
    G3_TEMP(2*I) <= G2_TEMP(2*I);
  END GENERATE EVEN_NODES_S3;
  
  -- NODE 5,7,9....63
  ODD_NODES_S3: FOR I IN 2 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S3_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G2_TEMP((2*I)+1),
	Pi => P2_TEMP((2*I)+1),
	Gj => G2_TEMP((2*I)-3),
	Pj => P2_TEMP((2*I)-3),
	P  => P3_TEMP((2*I)+1),
	G  => G3_TEMP((2*I)+1)
      );
   END GENERATE ODD_NODES_S3;

  -- STAGE 4
  -- NODE 0,1,2....8
  STAGE_4_INIT: FOR I IN 0 TO 8 GENERATE
    P4_TEMP(I) <= P3_TEMP(I);
    G4_TEMP(I) <= G3_TEMP(I);
  END GENERATE STAGE_4_INIT;

  -- NODE 10,12....62
  EVEN_NODES_S4: FOR I IN 5 TO (INPUT_WIDTH/2)-1 GENERATE
    P4_TEMP(2*I) <= P3_TEMP(2*I);
    G4_TEMP(2*I) <= G3_TEMP(2*I);
  END GENERATE EVEN_NODES_S4;

  -- NODE 9,11,....63
  ODD_NODES_S4: FOR I IN 4 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S4_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G3_TEMP((2*I)+1),
	Pi => P3_TEMP((2*I)+1),
	Gj => G3_TEMP((2*I)-7),
	Pj => P3_TEMP((2*I)-7),
	P  => P4_TEMP((2*I)+1),
	G  => G4_TEMP((2*I)+1)
      );
   END GENERATE ODD_NODES_S4;

  -- STAGE 5
  -- NODE 0,1,2....16
  STAGE_5_INIT: FOR I IN 0 TO 16 GENERATE
    P5_TEMP(I) <= P4_TEMP(I);
    G5_TEMP(I) <= G4_TEMP(I);
  END GENERATE STAGE_5_INIT;

  -- NODE 18,20....62
  EVEN_NODES_S5: FOR I IN 9 TO (INPUT_WIDTH/2)-1 GENERATE
    P5_TEMP(2*I) <= P4_TEMP(2*I);
    G5_TEMP(2*I) <= G4_TEMP(2*I);
  END GENERATE EVEN_NODES_S5;

  -- NODE 17,19....63
  ODD_NODES_S5: FOR I IN 8 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S5_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G4_TEMP((2*I)+1),
	Pi => P4_TEMP((2*I)+1),
	Gj => G4_TEMP((2*I)-15),
	Pj => P4_TEMP((2*I)-15),
	P  => P5_TEMP((2*I)+1),
	G  => G5_TEMP((2*I)+1)
      );
   END GENERATE ODD_NODES_S5;

  -- STAGE 6
  -- NODE 0,1,2....32
  STAGE_6_INIT: FOR I IN 0 TO 32 GENERATE
    P6_TEMP(I) <= P5_TEMP(I);
    G6_TEMP(I) <= G5_TEMP(I);
  END GENERATE STAGE_6_INIT;

  -- NODE 34,36....62
  EVEN_NODES_S6: FOR I IN 17 TO (INPUT_WIDTH/2)-1 GENERATE
    P6_TEMP(2*I) <= P5_TEMP(2*I);
    G6_TEMP(2*I) <= G5_TEMP(2*I);
  END GENERATE EVEN_NODES_S6;

  -- NODE 33,35....63
  ODD_NODES_S6: FOR I IN 16 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S6_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G5_TEMP((2*I)+1),
	Pi => P5_TEMP((2*I)+1),
	Gj => G5_TEMP((2*I)-31),
	Pj => P5_TEMP((2*I)-31),
	P  => P6_TEMP((2*I)+1),
	G  => G6_TEMP((2*I)+1)
      );
   END GENERATE ODD_NODES_S6;

  -- STAGE 7 (ADDITIONAL STAGE FOR HAN CARLSON ADDER)
  STAGE_7_INIT: FOR I IN 0 TO 1 GENERATE
    P7_TEMP(I) <= P6_TEMP(I);
    G7_TEMP(I) <= G6_TEMP(I);
  END GENERATE STAGE_7_INIT;

  -- NODE 2,4,6....62
  EVEN_NODES_S7: FOR I IN 1 TO (INPUT_WIDTH/2)-1 GENERATE
    PE_S7_I: PROCESS_ELEMENT PORT MAP
      (
	Gi => G6_TEMP(2*I),
	Pi => P6_TEMP(2*I),
	Gj => G6_TEMP((2*I)-1),
	Pj => P6_TEMP((2*I)-1),
	P  => P7_TEMP(2*I),
	G  => G7_TEMP(2*I)
      );
   END GENERATE EVEN_NODES_S7;

  -- NODE 3,5,7....63
  ODD_NODES_S7: FOR I IN 1 TO (INPUT_WIDTH/2)-1 GENERATE
    P7_TEMP((2*I)+1) <= P6_TEMP((2*I)+1);
    G7_TEMP((2*I)+1) <= G6_TEMP((2*I)+1);
  END GENERATE ODD_NODES_S7;

  -- POST PROCESSING: CALCULATING SUM
  S_TEMP(0) <= P0_TEMP(0);
  POST_PROCESSING: FOR I IN 1 TO INPUT_WIDTH-1 GENERATE
    S_TEMP(I) <= P0_TEMP(I) XOR G7_TEMP(I-1);
  END GENERATE POST_PROCESSING;

  S <= S_TEMP;
END BEHAVIORAL;  

