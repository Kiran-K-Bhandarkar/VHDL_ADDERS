-- IMPLEMENTED ADDER IS USING KOGGE STONE LOGIC

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY KS_ADDER IS 
GENERIC
(
  INPUT_WIDTH: INTEGER := 64
);

PORT
(
  NEG_B: IN STD_LOGIC;
  A, B: IN STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0);
  S: OUT STD_LOGIC_VECTOR(INPUT_WIDTH-1 DOWNTO 0)
);
END ENTITY KS_ADDER;

ARCHITECTURE BEHAVIORAL OF KS_ADDER IS

SIGNAL A_TEMP, B_TEMP, S_TEMP, 
P0_TEMP, G0_TEMP, P1_TEMP, G1_TEMP, 
P2_TEMP, G2_TEMP, P3_TEMP, G3_TEMP, 
P4_TEMP, G4_TEMP, P5_TEMP, G5_TEMP, 
P6_TEMP, G6_TEMP: STD_LOGIC_VECTOR(INPUT_WIDTH -1 DOWNTO 0) := (OTHERS => '0');

COMPONENT HALF_ADDER PORT
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END COMPONENT;

COMPONENT PROCESS_ELEMENT PORT
(
  Gi, Gj, Pi, Pj: IN STD_LOGIC;
  P, G: OUT STD_LOGIC
);
END COMPONENT;

BEGIN
  NEGATE_B: PROCESS(ALL)
    BEGIN
      IF NEG_B = '1' THEN
        B_TEMP <= NOT(B);
      ELSE
	B_TEMP <= B;
      END IF;
    END PROCESS;

  A_TEMP <= A;

  -- STAGE 0: OUTPUT FROM THE HALF ADDERS - PREPOCESSING STAGE
  PRE_PROCESSING: FOR I IN 0 TO INPUT_WIDTH-1 GENERATE
    HA_I: HALF_ADDER PORT MAP 
	(
	  A => A_TEMP(I), B => B_TEMP(I), 
	  S => P0_TEMP(I), C => G0_TEMP(I)
	);
  END GENERATE PRE_PROCESSING;
  
  -- STAGE 1
  P1_TEMP(0) <= P0_TEMP(0);
  G1_TEMP(0) <= G0_TEMP(0);

  STAGE_1: FOR I IN 1 TO INPUT_WIDTH-1 GENERATE
    PE_S1_I: PROCESS_ELEMENT PORT MAP
	(
	  Gi => G0_TEMP(I),
	  Pi => P0_TEMP(I),
	  Gj => G0_TEMP(I-1),
	  Pj => P0_TEMP(I-1),
	  P  => P1_TEMP(I),
	  G  => G1_TEMP(I)
	);
  END GENERATE STAGE_1;

  -- STAGE 2
  STAGE_2_INIT: FOR I IN 0 TO 1 GENERATE
    P2_TEMP(I) <= P1_TEMP(I);
    G2_TEMP(I) <= G1_TEMP(I);
  END GENERATE STAGE_2_INIT;

  STAGE_2: FOR I IN 2 TO INPUT_WIDTH-1 GENERATE
    PE_S2_I: PROCESS_ELEMENT PORT MAP
	(
	  Gi => G1_TEMP(I),
	  Pi => P1_TEMP(I),
	  Gj => G1_TEMP(I-2),
	  Pj => P1_TEMP(I-2),
	  P  => P2_TEMP(I),
	  G  => G2_TEMP(I)
	);
  END GENERATE STAGE_2;

  -- STAGE 3
  STAGE_3_INIT: FOR I IN 0 TO 3 GENERATE
    P3_TEMP(I) <= P2_TEMP(I);
    G3_TEMP(I) <= G2_TEMP(I);
  END GENERATE STAGE_3_INIT;

  STAGE_3: FOR I IN 4 TO INPUT_WIDTH-1 GENERATE
    PE_S3_I: PROCESS_ELEMENT PORT MAP
	(
	  Gi => G2_TEMP(I),
	  Pi => P2_TEMP(I),
	  Gj => G2_TEMP(I-4),
	  Pj => P2_TEMP(I-4),
	  P  => P3_TEMP(I),
	  G  => G3_TEMP(I)
	);
  END GENERATE STAGE_3;

  -- STAGE 4
  STAGE_4_INIT: FOR I IN 0 TO 7 GENERATE
    P4_TEMP(I) <= P3_TEMP(I);
    G4_TEMP(I) <= G3_TEMP(I);
  END GENERATE STAGE_4_INIT;

  STAGE_4: FOR I IN 8 TO INPUT_WIDTH-1 GENERATE
    PE_S4_I: PROCESS_ELEMENT PORT MAP
	(
	  Gi => G3_TEMP(I),
	  Pi => P3_TEMP(I),
	  Gj => G3_TEMP(I-8),
	  Pj => P3_TEMP(I-8),
	  P  => P4_TEMP(I),
	  G  => G4_TEMP(I)
	);
  END GENERATE STAGE_4;

  -- STAGE 5
  STAGE_5_INIT: FOR I IN 0 TO 15 GENERATE
    P5_TEMP(I) <= P4_TEMP(I);
    G5_TEMP(I) <= G4_TEMP(I);
  END GENERATE STAGE_5_INIT;

  STAGE_5: FOR I IN 16 TO INPUT_WIDTH-1 GENERATE
    PE_S5_I: PROCESS_ELEMENT PORT MAP
	(
	  Gi => G4_TEMP(I),
	  Pi => P4_TEMP(I),
	  Gj => G4_TEMP(I-16),
	  Pj => P4_TEMP(I-16),
	  P  => P5_TEMP(I),
	  G  => G5_TEMP(I)
	);
  END GENERATE STAGE_5;

  -- STAGE 6
  STAGE_6_INIT: FOR I IN 0 TO 31 GENERATE
    P6_TEMP(I) <= P5_TEMP(I);
    G6_TEMP(I) <= G5_TEMP(I);
  END GENERATE STAGE_6_INIT;

  STAGE_6: FOR I IN 32 TO INPUT_WIDTH-1 GENERATE
    PE_S6_I: PROCESS_ELEMENT PORT MAP
	(
	  Gi => G5_TEMP(I),
	  Pi => P5_TEMP(I),
	  Gj => G5_TEMP(I-32),
	  Pj => P5_TEMP(I-32),
	  P  => P6_TEMP(I),
	  G  => G6_TEMP(I)
	);
  END GENERATE STAGE_6;

  -- POST PROCESSING: CALCULATING SUM
  S_TEMP(0) <= P0_TEMP(0);
  POST_PROCESSING: FOR I IN 1 TO INPUT_WIDTH-1 GENERATE
    S_TEMP(I) <= P0_TEMP(I) XOR G6_TEMP(I-1);
  END GENERATE POST_PROCESSING;

  S <= S_TEMP;
END BEHAVIORAL;

