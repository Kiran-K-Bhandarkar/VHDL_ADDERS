LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CLA_64BIT IS PORT
(
  CI  : IN STD_LOGIC; 
  A, B: IN STD_LOGIC_VECTOR(63 DOWNTO 0);
  SUM : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END ENTITY CLA_64BIT;

ARCHITECTURE BEHAVIORAL OF CLA_64BIT IS
SIGNAL A_TEMP, B_TEMP, S_TEMP: STD_LOGIC_VECTOR(63 DOWNTO 0);
SIGNAL C_TEMP: STD_LOGIC_VECTOR(4 DOWNTO 0);

COMPONENT CLA_16BIT PORT
(
  A, B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
  CI   : IN STD_LOGIC;
  S    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
  CO   : OUT STD_LOGIC
);
END COMPONENT;

BEGIN
  A_TEMP    <= A;
  B_TEMP    <= B;
  C_TEMP(0) <= CI;

  -- 4x 16 BIT CLA CASCADED
  CLA_16B_0: CLA_16BIT PORT MAP
    (
      A  => A_TEMP(15 DOWNTO 0),
      B  => B_TEMP(15 DOWNTO 0),
      CI => C_TEMP(0),
      CO => C_TEMP(1),
      S  => S_TEMP(15 DOWNTO 0)
    );

  CLA_16B_1: CLA_16BIT PORT MAP
    (
      A  => A_TEMP(31 DOWNTO 16),
      B  => B_TEMP(31 DOWNTO 16),
      CI => C_TEMP(1),
      CO => C_TEMP(2),
      S  => S_TEMP(31 DOWNTO 16)
    );

  CLA_16B_2: CLA_16BIT PORT MAP
    (
      A  => A_TEMP(47 DOWNTO 32),
      B  => B_TEMP(47 DOWNTO 32),
      CI => C_TEMP(2),
      CO => C_TEMP(3),
      S  => S_TEMP(47 DOWNTO 32)
    );

  CLA_16B_3: CLA_16BIT PORT MAP
    (
      A  => A_TEMP(63 DOWNTO 48),
      B  => B_TEMP(63 DOWNTO 48),
      CI => C_TEMP(3),
      CO => C_TEMP(4),
      S  => S_TEMP(63 DOWNTO 48)
    );
  
  -- ASSIGNING OUTPUTS
  SUM  <= S_TEMP;
END BEHAVIORAL;