LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CLA_4BIT IS PORT
(
  A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
  CI   : IN STD_LOGIC;
  CO   : OUT STD_LOGIC;
  S    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END ENTITY CLA_4BIT;

ARCHITECTURE BEHAVIORAL OF CLA_4BIT IS 
SIGNAL A_TEMP, B_TEMP, G_PREPROCESS, P_PREPROCESS, S_TEMP: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL C_TEMP: STD_LOGIC_VECTOR(4 DOWNTO 0);

COMPONENT HALF_ADDER PORT
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END COMPONENT;

BEGIN
  A_TEMP    <= A;
  B_TEMP    <= B;
  C_TEMP(0) <= CI;

  -- PREPORCESSING STAGE: Pi AND Gi COMPUTING USING HALF ADDERS
  PREPROCESS: FOR I IN 0 TO 3 GENERATE
    HA_I: HALF_ADDER PORT MAP
      (
	A => A_TEMP(I),
	B => B_TEMP(I),
	S => P_PREPROCESS(I),
	C => G_PREPROCESS(I)
      );
    END GENERATE PREPROCESS;

  -- CARRY LOOK AHEAD BLOCK USING PREPOSSING ELEMENT
  CLA: FOR I IN 1 TO 4 GENERATE
    C_TEMP(I) <= G_PREPROCESS(I-1) OR (C_TEMP(I-1) AND P_PREPROCESS(I-1));
    END GENERATE CLA ;

  -- POST PROCESSING BLOCK
  POST_PROCESS: FOR I IN 0 TO 3 GENERATE
    S_TEMP(I) <= P_PREPROCESS(I) XOR C_TEMP(I);
  END GENERATE POST_PROCESS;

  -- ASSIGNING OUTPUT
  S  <= S_TEMP;
  CO <= C_TEMP(4);

END BEHAVIORAL;
	
	

