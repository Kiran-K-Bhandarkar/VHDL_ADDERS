LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FULL_ADDER IS PORT
(
  A,B,CI: IN STD_LOGIC;
  S, CO: OUT STD_LOGIC
);
END ENTITY FULL_ADDER;

ARCHITECTURE BEHAVIORAL OF FULL_ADDER IS
BEGIN
   S  <= A XOR B XOR CI;
   CO <= (A AND B) OR (CI AND (A XOR B));
END BEHAVIORAL;
