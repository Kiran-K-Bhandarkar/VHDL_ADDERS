LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RIPPLE_CARRY_ADDER IS PORT
(
  A,B  : IN STD_LOGIC_VECTOR(62 DOWNTO 0);
  CARRY: OUT STD_LOGIC;
  S    : OUT STD_LOGIC_VECTOR(62 DOWNTO 0)
);
END ENTITY RIPPLE_CARRY_ADDER;

ARCHITECTURE BEHAVIORAL OF RIPPLE_CARRY_ADDER IS
SIGNAL A_TEMP, B_TEMP, C_TEMP, S_TEMP: STD_LOGIC_VECTOR(62 DOWNTO 0) := (others => '0');

COMPONENT FULL_ADDER PORT
(
  A,B,CI: IN STD_LOGIC;
  S, CO: OUT STD_LOGIC
);
END COMPONENT;

COMPONENT HALF_ADDER PORT
(
  A, B: IN STD_LOGIC;
  S, C: OUT STD_LOGIC
);
END COMPONENT;
 
BEGIN
  A_TEMP <= A;
  B_TEMP <= B;

  -- LOWEST BITS USE HALF ADDER
  HA: HALF_ADDER PORT MAP
    (A => A_TEMP(0), B => B_TEMP(0), S => S_TEMP(0), C => C_TEMP(0));
  
  CARRY_CHAIN: FOR I IN 1 TO 62 GENERATE
    FA_I: FULL_ADDER PORT MAP
      (
	A  => A_TEMP(I),
	B  => B_TEMP(I),
	CI => C_TEMP(I-1),
	CO => C_TEMP(I),
	S  => S_TEMP(I)
      );
    END GENERATE CARRY_CHAIN;

  -- OUTPUT CONCATINATING THE SUM AND THE CARRY BIT OF THE LAST FULL ADDER
  S     <= S_TEMP;
  CARRY <= C_TEMP(62);
END BEHAVIORAL;
