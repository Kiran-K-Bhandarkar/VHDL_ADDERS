LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CLA_16BIT IS PORT
(
  A, B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
  CI   : IN STD_LOGIC;
  S    : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
  CO   : OUT STD_LOGIC
);
END ENTITY CLA_16BIT;

ARCHITECTURE BEHAVIORAL OF CLA_16BIT IS
SIGNAL A_TEMP, B_TEMP, S_TEMP: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL C_TEMP: STD_LOGIC_VECTOR(4 DOWNTO 0);

COMPONENT CLA_4BIT PORT
(
  A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
  CI   : IN STD_LOGIC;
  CO   : OUT STD_LOGIC;
  S    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);
END COMPONENT; 

BEGIN
  A_TEMP    <= A;
  B_TEMP    <= B;
  C_TEMP(0) <= CI;

  -- 4x 4 BIT CLA CASCADED
  CLA_4B_0: CLA_4BIT PORT MAP
    (
      A  => A_TEMP(3 DOWNTO 0),
      B  => B_TEMP(3 DOWNTO 0),
      CI => C_TEMP(0),
      CO => C_TEMP(1),
      S  => S_TEMP(3 DOWNTO 0)
    );

  CLA_4B_1: CLA_4BIT PORT MAP
    (
      A  => A_TEMP(7 DOWNTO 4),
      B  => B_TEMP(7 DOWNTO 4),
      CI => C_TEMP(1),
      CO => C_TEMP(2),
      S  => S_TEMP(7 DOWNTO 4)
    );

  CLA_4B_2: CLA_4BIT PORT MAP
    (
      A  => A_TEMP(11 DOWNTO 8),
      B  => B_TEMP(11 DOWNTO 8),
      CI => C_TEMP(2),
      CO => C_TEMP(3),
      S  => S_TEMP(11 DOWNTO 8)
    );

  CLA_4B_3: CLA_4BIT PORT MAP
    (
      A  => A_TEMP(15 DOWNTO 12),
      B  => B_TEMP(15 DOWNTO 12),
      CI => C_TEMP(3),
      CO => C_TEMP(4),
      S  => S_TEMP(15 DOWNTO 12)
    );

  -- ASSIGNING OUTPUTS
  S  <= S_TEMP;
  CO <= C_TEMP(4);

END BEHAVIORAL;